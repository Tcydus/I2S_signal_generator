library verilog;
use verilog.vl_types.all;
entity DAC_Input_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        RST_BTN         : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end DAC_Input_vlg_sample_tst;
