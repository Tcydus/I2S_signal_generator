library verilog;
use verilog.vl_types.all;
entity DAC_Input_vlg_vec_tst is
end DAC_Input_vlg_vec_tst;
